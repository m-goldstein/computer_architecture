
import sourcemux::*;
import validmux::*;
import datamux::*;
import dirtymux::*;
import waymux::*;
import tagmux::*;
import destmux::*;
import waymux::*;
import tagmux::*;
import hitmux::*;

